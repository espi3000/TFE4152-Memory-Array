*************************************
* 3 INPUT NAND GATE
*************************************
.subckt 3_in_nand y a b c vdd vss
.include param.cir
xmp1 y a vdd vdd pmos1v l=lp w=wp
xmp2 y b vdd vdd pmos1v l=lp w=wp
xmp3 y c vdd vdd pmos1v l=lp w=wp
xmn1 y a 1 1 nmos1v l=ln w=wn
xmn2 1 b 2 2 nmos1v l=ln w=wn
xmn3 2 c vss vss nmos1v l=ln w=wn
.ends

*************************************
* 2 INPUT NAND GATE
*************************************
.subckt 2_in_nand y a b vdd vss
.include param.cir
xmp1 y a vdd vdd pmos1v l=lp w=wp
xmp2 y b vdd vdd pmos1v l=lp w=wp
xmn1 y a 1 1 nmos1v l=ln w=wn
xmn2 1 b vss vss nmos1v l=ln w=wn
.ends
*************************************
* PARAMS
*************************************
.param ln = 150n
.param lp = 150n
.param wn = 150n
.param wp = 1500n
.param vh = 0.45

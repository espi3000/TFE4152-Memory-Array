*************************************
* PARAMS
*************************************
.param ln = 0.1u
.param lp = 0.1u
.param wn = 0.1u
.param wp = 0.1u

*************************************
* PARAMS
*************************************
.param ln = 90n
.param lp = 90n
.param wn = 90n
.param wp = 300n

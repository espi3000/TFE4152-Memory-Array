* 3 INPUT NOR GATE
.subckt 3_in_nor y a b c vdd vss
.include param.cir
xmp1 1 a vdd vdd pmos1v l=lp w=wp
xmp2 2 b 1 1 pmos1v l=lp w=wp
xmp3 y c 2 2 pmos1v l=lp w=wp
xmn1 y a vss vss pmos1v l=lp w=wp
xmn2 y b vss vss pmos1v l=lp w=wp
xmn3 y c vss vss pmos1v l=lp w=wp
.ends

* 2 INPUT NOR GATE
.subckt 2_in_nor y a b vdd vss
.include param.cir
xmp1 1 a vdd vdd pmos1v l=lp w=wp
xmp2 y b 1 1 pmos1v l=lp w=wp
xmn1 y a vss vss pmos1v l=lp w=wp
xmn2 y b vss vss pmos1v l=lp w=wp
.ends